VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_tpm2137
  CLASS BLOCK ;
  FOREIGN wrapped_tpm2137 ;
  ORIGIN 0.000 0.000 ;
  SIZE 130.000 BY 210.000 ;
  PIN active
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 201.320 130.000 201.920 ;
    END
  END active
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 57.160 130.000 57.760 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 206.000 7.730 210.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 4.000 110.800 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 206.000 115.370 210.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 206.000 92.370 210.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.800 4.000 124.400 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 206.000 40.850 210.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 0.000 37.170 4.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 187.720 130.000 188.320 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 15.000 130.000 15.600 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.490 206.000 110.770 210.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 4.000 138.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.560 4.000 180.160 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 97.960 130.000 98.560 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 186.360 4.000 186.960 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 206.000 59.250 210.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 194.520 130.000 195.120 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 1.400 130.000 2.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 70.760 130.000 71.360 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 206.000 54.650 210.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 111.560 130.000 112.160 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 4.000 117.600 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 0.000 50.970 4.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 28.600 130.000 29.200 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.000 4.000 151.600 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.970 206.000 36.250 210.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 77.560 130.000 78.160 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 118.360 130.000 118.960 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 206.000 68.450 210.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 91.160 130.000 91.760 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 206.000 73.050 210.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 206.000 83.170 210.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 206.000 101.570 210.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 206.000 129.170 210.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 174.120 130.000 174.720 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 4.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.650 206.000 16.930 210.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 0.000 61.090 4.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 4.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 180.920 130.000 181.520 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.530 0.000 121.810 4.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 140.120 130.000 140.720 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 206.000 50.050 210.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 4.000 97.200 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 206.000 27.050 210.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.570 206.000 63.850 210.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.810 0.000 107.090 4.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.490 0.000 41.770 4.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 63.960 130.000 64.560 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 206.000 31.650 210.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 146.920 130.000 147.520 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.290 0.000 9.570 4.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.130 0.000 126.410 4.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 50.360 130.000 50.960 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 206.000 124.570 210.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.960 4.000 166.560 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 0.000 112.610 4.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 0.000 56.490 4.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.800 4.000 158.400 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 160.520 130.000 161.120 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 4.000 90.400 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 21.800 130.000 22.400 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.960 4.000 200.560 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 206.000 12.330 210.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 4.000 131.200 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 0.000 97.890 4.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 0.000 14.170 4.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 4.000 83.600 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 8.200 130.000 8.800 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 125.160 130.000 125.760 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 84.360 130.000 84.960 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 4.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.200 4.000 144.800 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 42.200 130.000 42.800 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 4.000 104.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 153.720 130.000 154.320 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.930 0.000 117.210 4.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 167.320 130.000 167.920 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.010 0.000 70.290 4.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 0.000 88.690 4.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.850 206.000 3.130 210.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 206.000 45.450 210.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 206.000 87.770 210.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 0.000 23.370 4.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 0.000 4.970 4.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 206.000 106.170 210.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 206.000 78.570 210.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 0.000 65.690 4.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 206.000 119.970 210.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 35.400 130.000 36.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 4.000 193.760 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 4.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.090 0.000 46.370 4.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 133.320 130.000 133.920 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 4.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 206.000 96.970 210.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.760 4.000 207.360 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.170 206.000 22.450 210.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.010 0.000 93.290 4.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.760 4.000 173.360 ;
    END
  END io_out[9]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 24.545 10.640 26.145 198.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 64.195 10.640 65.795 198.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 103.850 10.640 105.450 198.800 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 44.370 10.640 45.970 198.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 84.025 10.640 85.625 198.800 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 104.760 130.000 105.360 ;
    END
  END wb_clk_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 125.435 198.645 ;
      LAYER met1 ;
        RECT 0.070 10.640 129.190 198.800 ;
      LAYER met2 ;
        RECT 0.100 205.720 2.570 207.245 ;
        RECT 3.410 205.720 7.170 207.245 ;
        RECT 8.010 205.720 11.770 207.245 ;
        RECT 12.610 205.720 16.370 207.245 ;
        RECT 17.210 205.720 21.890 207.245 ;
        RECT 22.730 205.720 26.490 207.245 ;
        RECT 27.330 205.720 31.090 207.245 ;
        RECT 31.930 205.720 35.690 207.245 ;
        RECT 36.530 205.720 40.290 207.245 ;
        RECT 41.130 205.720 44.890 207.245 ;
        RECT 45.730 205.720 49.490 207.245 ;
        RECT 50.330 205.720 54.090 207.245 ;
        RECT 54.930 205.720 58.690 207.245 ;
        RECT 59.530 205.720 63.290 207.245 ;
        RECT 64.130 205.720 67.890 207.245 ;
        RECT 68.730 205.720 72.490 207.245 ;
        RECT 73.330 205.720 78.010 207.245 ;
        RECT 78.850 205.720 82.610 207.245 ;
        RECT 83.450 205.720 87.210 207.245 ;
        RECT 88.050 205.720 91.810 207.245 ;
        RECT 92.650 205.720 96.410 207.245 ;
        RECT 97.250 205.720 101.010 207.245 ;
        RECT 101.850 205.720 105.610 207.245 ;
        RECT 106.450 205.720 110.210 207.245 ;
        RECT 111.050 205.720 114.810 207.245 ;
        RECT 115.650 205.720 119.410 207.245 ;
        RECT 120.250 205.720 124.010 207.245 ;
        RECT 124.850 205.720 128.610 207.245 ;
        RECT 0.100 4.280 129.160 205.720 ;
        RECT 0.650 3.670 4.410 4.280 ;
        RECT 5.250 3.670 9.010 4.280 ;
        RECT 9.850 3.670 13.610 4.280 ;
        RECT 14.450 3.670 18.210 4.280 ;
        RECT 19.050 3.670 22.810 4.280 ;
        RECT 23.650 3.670 27.410 4.280 ;
        RECT 28.250 3.670 32.010 4.280 ;
        RECT 32.850 3.670 36.610 4.280 ;
        RECT 37.450 3.670 41.210 4.280 ;
        RECT 42.050 3.670 45.810 4.280 ;
        RECT 46.650 3.670 50.410 4.280 ;
        RECT 51.250 3.670 55.930 4.280 ;
        RECT 56.770 3.670 60.530 4.280 ;
        RECT 61.370 3.670 65.130 4.280 ;
        RECT 65.970 3.670 69.730 4.280 ;
        RECT 70.570 3.670 74.330 4.280 ;
        RECT 75.170 3.670 78.930 4.280 ;
        RECT 79.770 3.670 83.530 4.280 ;
        RECT 84.370 3.670 88.130 4.280 ;
        RECT 88.970 3.670 92.730 4.280 ;
        RECT 93.570 3.670 97.330 4.280 ;
        RECT 98.170 3.670 101.930 4.280 ;
        RECT 102.770 3.670 106.530 4.280 ;
        RECT 107.370 3.670 112.050 4.280 ;
        RECT 112.890 3.670 116.650 4.280 ;
        RECT 117.490 3.670 121.250 4.280 ;
        RECT 122.090 3.670 125.850 4.280 ;
        RECT 126.690 3.670 129.160 4.280 ;
      LAYER met3 ;
        RECT 4.400 206.360 126.000 207.225 ;
        RECT 4.000 202.320 126.000 206.360 ;
        RECT 4.000 200.960 125.600 202.320 ;
        RECT 4.400 200.920 125.600 200.960 ;
        RECT 4.400 199.560 126.000 200.920 ;
        RECT 4.000 195.520 126.000 199.560 ;
        RECT 4.000 194.160 125.600 195.520 ;
        RECT 4.400 194.120 125.600 194.160 ;
        RECT 4.400 192.760 126.000 194.120 ;
        RECT 4.000 188.720 126.000 192.760 ;
        RECT 4.000 187.360 125.600 188.720 ;
        RECT 4.400 187.320 125.600 187.360 ;
        RECT 4.400 185.960 126.000 187.320 ;
        RECT 4.000 181.920 126.000 185.960 ;
        RECT 4.000 180.560 125.600 181.920 ;
        RECT 4.400 180.520 125.600 180.560 ;
        RECT 4.400 179.160 126.000 180.520 ;
        RECT 4.000 175.120 126.000 179.160 ;
        RECT 4.000 173.760 125.600 175.120 ;
        RECT 4.400 173.720 125.600 173.760 ;
        RECT 4.400 172.360 126.000 173.720 ;
        RECT 4.000 168.320 126.000 172.360 ;
        RECT 4.000 166.960 125.600 168.320 ;
        RECT 4.400 166.920 125.600 166.960 ;
        RECT 4.400 165.560 126.000 166.920 ;
        RECT 4.000 161.520 126.000 165.560 ;
        RECT 4.000 160.120 125.600 161.520 ;
        RECT 4.000 158.800 126.000 160.120 ;
        RECT 4.400 157.400 126.000 158.800 ;
        RECT 4.000 154.720 126.000 157.400 ;
        RECT 4.000 153.320 125.600 154.720 ;
        RECT 4.000 152.000 126.000 153.320 ;
        RECT 4.400 150.600 126.000 152.000 ;
        RECT 4.000 147.920 126.000 150.600 ;
        RECT 4.000 146.520 125.600 147.920 ;
        RECT 4.000 145.200 126.000 146.520 ;
        RECT 4.400 143.800 126.000 145.200 ;
        RECT 4.000 141.120 126.000 143.800 ;
        RECT 4.000 139.720 125.600 141.120 ;
        RECT 4.000 138.400 126.000 139.720 ;
        RECT 4.400 137.000 126.000 138.400 ;
        RECT 4.000 134.320 126.000 137.000 ;
        RECT 4.000 132.920 125.600 134.320 ;
        RECT 4.000 131.600 126.000 132.920 ;
        RECT 4.400 130.200 126.000 131.600 ;
        RECT 4.000 126.160 126.000 130.200 ;
        RECT 4.000 124.800 125.600 126.160 ;
        RECT 4.400 124.760 125.600 124.800 ;
        RECT 4.400 123.400 126.000 124.760 ;
        RECT 4.000 119.360 126.000 123.400 ;
        RECT 4.000 118.000 125.600 119.360 ;
        RECT 4.400 117.960 125.600 118.000 ;
        RECT 4.400 116.600 126.000 117.960 ;
        RECT 4.000 112.560 126.000 116.600 ;
        RECT 4.000 111.200 125.600 112.560 ;
        RECT 4.400 111.160 125.600 111.200 ;
        RECT 4.400 109.800 126.000 111.160 ;
        RECT 4.000 105.760 126.000 109.800 ;
        RECT 4.000 104.400 125.600 105.760 ;
        RECT 4.400 104.360 125.600 104.400 ;
        RECT 4.400 103.000 126.000 104.360 ;
        RECT 4.000 98.960 126.000 103.000 ;
        RECT 4.000 97.600 125.600 98.960 ;
        RECT 4.400 97.560 125.600 97.600 ;
        RECT 4.400 96.200 126.000 97.560 ;
        RECT 4.000 92.160 126.000 96.200 ;
        RECT 4.000 90.800 125.600 92.160 ;
        RECT 4.400 90.760 125.600 90.800 ;
        RECT 4.400 89.400 126.000 90.760 ;
        RECT 4.000 85.360 126.000 89.400 ;
        RECT 4.000 84.000 125.600 85.360 ;
        RECT 4.400 83.960 125.600 84.000 ;
        RECT 4.400 82.600 126.000 83.960 ;
        RECT 4.000 78.560 126.000 82.600 ;
        RECT 4.000 77.160 125.600 78.560 ;
        RECT 4.000 75.840 126.000 77.160 ;
        RECT 4.400 74.440 126.000 75.840 ;
        RECT 4.000 71.760 126.000 74.440 ;
        RECT 4.000 70.360 125.600 71.760 ;
        RECT 4.000 69.040 126.000 70.360 ;
        RECT 4.400 67.640 126.000 69.040 ;
        RECT 4.000 64.960 126.000 67.640 ;
        RECT 4.000 63.560 125.600 64.960 ;
        RECT 4.000 62.240 126.000 63.560 ;
        RECT 4.400 60.840 126.000 62.240 ;
        RECT 4.000 58.160 126.000 60.840 ;
        RECT 4.000 56.760 125.600 58.160 ;
        RECT 4.000 55.440 126.000 56.760 ;
        RECT 4.400 54.040 126.000 55.440 ;
        RECT 4.000 51.360 126.000 54.040 ;
        RECT 4.000 49.960 125.600 51.360 ;
        RECT 4.000 48.640 126.000 49.960 ;
        RECT 4.400 47.240 126.000 48.640 ;
        RECT 4.000 43.200 126.000 47.240 ;
        RECT 4.000 41.840 125.600 43.200 ;
        RECT 4.400 41.800 125.600 41.840 ;
        RECT 4.400 40.440 126.000 41.800 ;
        RECT 4.000 36.400 126.000 40.440 ;
        RECT 4.000 35.040 125.600 36.400 ;
        RECT 4.400 35.000 125.600 35.040 ;
        RECT 4.400 33.640 126.000 35.000 ;
        RECT 4.000 29.600 126.000 33.640 ;
        RECT 4.000 28.240 125.600 29.600 ;
        RECT 4.400 28.200 125.600 28.240 ;
        RECT 4.400 26.840 126.000 28.200 ;
        RECT 4.000 22.800 126.000 26.840 ;
        RECT 4.000 21.440 125.600 22.800 ;
        RECT 4.400 21.400 125.600 21.440 ;
        RECT 4.400 20.040 126.000 21.400 ;
        RECT 4.000 16.000 126.000 20.040 ;
        RECT 4.000 14.640 125.600 16.000 ;
        RECT 4.400 14.600 125.600 14.640 ;
        RECT 4.400 13.240 126.000 14.600 ;
        RECT 4.000 9.200 126.000 13.240 ;
        RECT 4.000 7.840 125.600 9.200 ;
        RECT 4.400 7.800 125.600 7.840 ;
        RECT 4.400 6.975 126.000 7.800 ;
  END
END wrapped_tpm2137
END LIBRARY

